library verilog;
use verilog.vl_types.all;
entity randnum_vlg_vec_tst is
end randnum_vlg_vec_tst;

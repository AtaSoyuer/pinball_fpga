module score (input wire i_clk,         // base clock
						input wire i_ani_stb,     // animation clock: pixel clock is 1 pix/frame
						input wire i_rst,         // reset: returns animation to starting position
						input wire i_animate,     // animate when input is high
						input [9:0] x, y,
						input [11:0] score,
						output reg a0,a1,a2,a3,a4,a5,a6,
						output reg b0,b1,b2,b3,b4,b5,b6,
						output reg c0,c1,c2,c3,c4,c5,c6
						
						 );




reg [3:0] A, B, C ;

initial
begin
A=0;
B=0;
C=0;

end


    

 integer i;
 always @(score)

 begin
 
 if(i_animate)
 begin
  // sets
  A = 4'd0;
  B = 4'd0;
  C = 4'd0;
  
  
  for(i=11 ; i>=0 ; i=i-1)
	begin
		if( A >= 5)
				A = A +3;
		if( B>= 5)
				B = B + 3;
		if( C >= 5)
				C = C +3;
	 
			// shifts
	   A = A << 1;
		A[0] = B[3];
		B = B << 1;
		C[0] = C[3];
		C = C << 1;
		C[0] = score[i] ;
	 end
 end
 end

						 
// Seven segment creation	
always @ (posedge i_clk)
begin
case (A)
0:
begin 
a0=((x>=10)&&(x<=35)&&(y==50));
a1=((y>=50)&&(y<=75)&&(x==35));
a2=((y>=75)&&(y<=100)&&(x==35));
a3=((x>=10)&&(x<=35)&&(y==100));
a4=((y>=75)&&(y<=100)&&(x==10));
a5=((y>=50)&&(y<=75)&&(x==10));
a6=0;
end
1:
begin 
a0=0;
a1=((y>=50)&&(y<=75)&&(x==35));
a2=((y>=75)&&(y<=100)&&(x==35));
a3=0;
a4=0;
a5=0;
a6=0;
end
2:
begin 
a0=((x>=10)&&(x<=35)&&(y==50));
a1=((y>=50)&&(y<=75)&&(x==35));
a2=0;
a3=((x>=10)&&(x<=35)&&(y==100));
a4=((y>=75)&&(y<=100)&&(x==10));
a5=0;
a6=((x>=10)&&(x<=35)&&(y==75));
end
3:
begin 
a0=((x>=10)&&(x<=35)&&(y==50));
a1=((y>=50)&&(y<=75)&&(x==35));
a2=((y>=75)&&(y<=100)&&(x==35));
a3=((x>=10)&&(x<=35)&&(y==100));
a4=0;
a5=0;
a6=((x>=10)&&(x<=35)&&(y==75));
end
4:
begin 
a0=0;
a1=((y>=50)&&(y<=75)&&(x==35));
a2=((y>=75)&&(y<=100)&&(x==35));
a3=0;
a4=0;
a5=((y>=50)&&(y<=75)&&(x==10));
a6=((x>=10)&&(x<=35)&&(y==75));
end
5:
begin 
a0=((x>=10)&&(x<=35)&&(y==50));
a1=0;
a2=((y>=75)&&(y<=100)&&(x==35));
a3=((x>=10)&&(x<=35)&&(y==100));
a4=0;
a5=((y>=50)&&(y<=75)&&(x==10));
a6=((x>=10)&&(x<=35)&&(y==75));
end
6:
begin 
a0=((x>=10)&&(x<=35)&&(y==50));
a1=0;
a2=((y>=75)&&(y<=100)&&(x==35));
a3=((x>=10)&&(x<=35)&&(y==100));
a4=((y>=75)&&(y<=100)&&(x==10));
a5=((y>=50)&&(y<=75)&&(x==10));
a6=((x>=10)&&(x<=35)&&(y==75));
end
7:
begin 
a0=((x>=10)&&(x<=35)&&(y==50));
a1=((y>=50)&&(y<=75)&&(x==35));
a2=((y>=75)&&(y<=100)&&(x==35));
a3=0;
a4=0;
a5=0;
a6=0;
end
8:
begin 
a0=((x>=10)&&(x<=35)&&(y==50));
a1=((y>=50)&&(y<=75)&&(x==35));
a2=((y>=75)&&(y<=100)&&(x==35));
a3=((x>=10)&&(x<=35)&&(y==100));
a4=((y>=75)&&(y<=100)&&(x==10));
a5=((y>=50)&&(y<=75)&&(x==10));
a6=((x>=10)&&(x<=35)&&(y==75));
end
9:
begin 
a0=((x>=10)&&(x<=35)&&(y==50));
a1=((y>=50)&&(y<=75)&&(x==35));
a2=((y>=75)&&(y<=100)&&(x==35));
a3=((x>=10)&&(x<=35)&&(y==100));
a4=0;
a5=((y>=50)&&(y<=75)&&(x==10));
a6=((x>=10)&&(x<=35)&&(y==75));
end
endcase
end


						 
always @ (posedge i_clk)
begin


case (B)
0:
begin 
b0=((x>=45)&&(x<=70)&&(y==50));
b1=((y>=50)&&(y<=75)&&(x==70));
b2=((y>=75)&&(y<=100)&&(x==70));
b3=((x>=45)&&(x<=70)&&(y==100));
b4=((y>=75)&&(y<=100)&&(x==45));
b5=((y>=50)&&(y<=75)&&(x==45));
b6=0;
end
1:
begin 
b0=0;
b1=((y>=50)&&(y<=75)&&(x==70));
b2=((y>=75)&&(y<=100)&&(x==70));
b3=0;
b4=0;
b5=0;
b6=0;
end
2:
begin 
b0=((x>=45)&&(x<=70)&&(y==50));
b1=((y>=50)&&(y<=75)&&(x==70));
b2=0;
b3=((x>=45)&&(x<=70)&&(y==100));
b4=((y>=75)&&(y<=100)&&(x==45));
b5=0;
b6=((x>=45)&&(x<=70)&&(y==75));
end
3:
begin 
b0=((x>=45)&&(x<=70)&&(y==50));
b1=((y>=50)&&(y<=75)&&(x==70));
b2=((y>=75)&&(y<=100)&&(x==70));
b3=((x>=45)&&(x<=70)&&(y==100));
b4=0;
b5=0;
b6=((x>=45)&&(x<=70)&&(y==75));
end
4:
begin 
b0=0;
b1=((y>=50)&&(y<=75)&&(x==70));
b2=((y>=75)&&(y<=100)&&(x==70));
b3=0;
b4=0;
b5=((y>=50)&&(y<=75)&&(x==45));
b6=((x>=45)&&(x<=70)&&(y==75));
end
5:
begin 
b0=((x>=45)&&(x<=70)&&(y==50));
b1=0;
b2=((y>=75)&&(y<=100)&&(x==70));
b3=((x>=45)&&(x<=70)&&(y==100));
b4=0;
b5=((y>=50)&&(y<=75)&&(x==45));
b6=((x>=45)&&(x<=70)&&(y==75));
end
6:
begin 
b0=((x>=45)&&(x<=70)&&(y==50));
b1=0;
b2=((y>=75)&&(y<=100)&&(x==70));
b3=((x>=45)&&(x<=70)&&(y==100));
b4=((y>=75)&&(y<=100)&&(x==45));
b5=((y>=50)&&(y<=75)&&(x==45));
b6=((x>=45)&&(x<=70)&&(y==75));
end
7:
begin 
b0=((x>=45)&&(x<=70)&&(y==50));
b1=((y>=50)&&(y<=75)&&(x==70));
b2=((y>=75)&&(y<=100)&&(x==70));
b3=0;
b4=0;
b5=0;
b6=0;
end
8:
begin 
b0=((x>=45)&&(x<=70)&&(y==50));
b1=((y>=50)&&(y<=75)&&(x==70));
b2=((y>=75)&&(y<=100)&&(x==70));
b3=((x>=45)&&(x<=70)&&(y==100));
b4=((y>=75)&&(y<=100)&&(x==45));
b5=((y>=50)&&(y<=75)&&(x==45));
b6=((x>=45)&&(x<=70)&&(y==75));
end
9:
begin 
b0=((x>=45)&&(x<=70)&&(y==50));
b1=((y>=50)&&(y<=75)&&(x==70));
b2=((y>=75)&&(y<=100)&&(x==70));
b3=((x>=45)&&(x<=70)&&(y==100));
b4=0;
b5=((y>=50)&&(y<=75)&&(x==45));
b6=((x>=45)&&(x<=70)&&(y==75));
end
endcase
end



always @ (posedge i_clk)
begin

case (C)
0:
begin 
c0=((x>=80)&&(x<=105)&&(y==50));
c1=((y>=50)&&(y<=75)&&(x==105));
c2=((y>=75)&&(y<=100)&&(x==105));
c3=((x>=80)&&(x<=105)&&(y==100));
c4=((y>=75)&&(y<=100)&&(x==80));
c5=((y>=50)&&(y<=75)&&(x==80));
c6=0;
end
1:
begin 
c0=0;
c1=((y>=50)&&(y<=75)&&(x==105));
c2=((y>=75)&&(y<=100)&&(x==105));
c3=0;
c4=0;
c5=0;
c6=0;
end
2:
begin 
c0=((x>=80)&&(x<=105)&&(y==50));
c1=((y>=50)&&(y<=75)&&(x==105));
c2=0;
c3=((x>=80)&&(x<=105)&&(y==100));
c4=((y>=75)&&(y<=100)&&(x==80));
c5=0;
c6=((x>=80)&&(x<=105)&&(y==75));
end
3:
begin 
c0=((x>=80)&&(x<=105)&&(y==50));
c1=((y>=50)&&(y<=75)&&(x==105));
c2=((y>=75)&&(y<=100)&&(x==105));
c3=((x>=80)&&(x<=105)&&(y==100));
c4=0;
c5=0;
c6=((x>=80)&&(x<=105)&&(y==75));
end
4:
begin 
c0=0;
c1=((y>=50)&&(y<=75)&&(x==105));
c2=((y>=75)&&(y<=100)&&(x==105));
c3=0;
c4=0;
c5=((y>=50)&&(y<=75)&&(x==80));
c6=((x>=80)&&(x<=105)&&(y==75));
end
5:
begin 
c0=((x>=80)&&(x<=105)&&(y==50));
c1=0;
c2=((y>=75)&&(y<=100)&&(x==105));
c3=((x>=80)&&(x<=105)&&(y==100));
c4=0;
c5=((y>=50)&&(y<=75)&&(x==80));
c6=((x>=80)&&(x<=105)&&(y==75));
end
6:
begin 
c0=0;
c1=((y>=50)&&(y<=75)&&(x==105));
c2=((y>=75)&&(y<=100)&&(x==105));
c3=((x>=80)&&(x<=105)&&(y==100));
c4=((y>=75)&&(y<=100)&&(x==80));
c5=((y>=50)&&(y<=75)&&(x==80));
c6=((x>=80)&&(x<=105)&&(y==75));
end
7:
begin 
c0=((x>=80)&&(x<=105)&&(y==50));
c1=((y>=50)&&(y<=75)&&(x==105));
c2=((y>=75)&&(y<=100)&&(x==105));
c3=0;
c4=0;
c5=0;
c6=0;
end
8:
begin 
c0=((x>=80)&&(x<=105)&&(y==50));
c1=((y>=50)&&(y<=75)&&(x==105));
c2=((y>=75)&&(y<=100)&&(x==105));
c3=((x>=80)&&(x<=105)&&(y==100));
c4=((y>=75)&&(y<=100)&&(x==80));
c5=((y>=50)&&(y<=75)&&(x==80));
c6=((x>=80)&&(x<=105)&&(y==75));
end
9:
begin 
c0=((x>=80)&&(x<=105)&&(y==50));
c1=((y>=50)&&(y<=75)&&(x==105));
c2=((y>=75)&&(y<=100)&&(x==105));
c3=((x>=80)&&(x<=105)&&(y==100));
c4=0;
c5=((y>=50)&&(y<=75)&&(x==80));
c6=((x>=80)&&(x<=105)&&(y==75));
end
endcase
end					 
endmodule						 
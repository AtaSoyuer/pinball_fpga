library verilog;
use verilog.vl_types.all;
entity clk_en_vlg_vec_tst is
end clk_en_vlg_vec_tst;

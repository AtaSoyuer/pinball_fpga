library verilog;
use verilog.vl_types.all;
entity hexagon_vlg_vec_tst is
end hexagon_vlg_vec_tst;

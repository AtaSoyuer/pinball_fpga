library verilog;
use verilog.vl_types.all;
entity hexagon_vlg_check_tst is
    port(
        hexagon         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end hexagon_vlg_check_tst;
